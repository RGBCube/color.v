module color

pub type Color = BasicColor | TrueColor
