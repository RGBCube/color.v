module main

import color

fn main() {
	println(color.red.color('Hello World'))
	println(color.bold.color('Hello World'))
}
