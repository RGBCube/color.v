module main

import color

fn main() {
	color.red.cprintln('Hello World')
	color.bold.cprintln('Hello World')
}
