module main

import color

fn main() {
	println(color.red.apply('Hello World'))
	println(color.bold.apply('Hello World'))
}
